`define N 9		/* для хранения количества роутеров и эмуряции пакета */
`define N2 17   /* это размер входящего и выходящего пакетов - 1 бит для эмуляции и K*2 бит для передачи двух чисел (шагов по первой и по второй образующим)*/
`define N_COUNT 144  /* это количество роутеров с отсчетом с нулевого, поэтому это значение всегда будет на один меньше от счетного количества*/

module toplevel_apo_144_nodes(
	clk,

	sw_on,
	sw_sel_data,
	sw_sel_router,
	key_inc,
	key_dec,

	out_data,

	hex_data,
	hex_router
);
	input clk;

	input sw_on;
	input sw_sel_data;
	input sw_sel_router;
	input key_inc;
	input key_dec;

	output wire[143:0] out_data;
	output wire[6:0] hex_data;
	output wire[6:0] hex_router;

	wire[`N2-1:0] out_router1;
	wire[`N2-1:0] out_router2;
	wire[`N2-1:0] out_router3;
	wire[`N2-1:0] out_router4;
	wire[`N2-1:0] out_router5;
	wire[`N2-1:0] out_router6;
	wire[`N2-1:0] out_router7;
	wire[`N2-1:0] out_router8;
	wire[`N2-1:0] out_router9;
	wire[`N2-1:0] out_router10;
	wire[`N2-1:0] out_router11;
	wire[`N2-1:0] out_router12;
	wire[`N2-1:0] out_router13;
	wire[`N2-1:0] out_router14;
	wire[`N2-1:0] out_router15;
	wire[`N2-1:0] out_router16;
	wire[`N2-1:0] out_router17;
	wire[`N2-1:0] out_router18;
	wire[`N2-1:0] out_router19;
	wire[`N2-1:0] out_router20;
	wire[`N2-1:0] out_router21;
	wire[`N2-1:0] out_router22;
	wire[`N2-1:0] out_router23;
	wire[`N2-1:0] out_router24;
	wire[`N2-1:0] out_router25;
	wire[`N2-1:0] out_router26;
	wire[`N2-1:0] out_router27;
	wire[`N2-1:0] out_router28;
	wire[`N2-1:0] out_router29;
	wire[`N2-1:0] out_router30;
	wire[`N2-1:0] out_router31;
	wire[`N2-1:0] out_router32;
	wire[`N2-1:0] out_router33;
	wire[`N2-1:0] out_router34;
	wire[`N2-1:0] out_router35;
	wire[`N2-1:0] out_router36;
	wire[`N2-1:0] out_router37;
	wire[`N2-1:0] out_router38;
	wire[`N2-1:0] out_router39;
	wire[`N2-1:0] out_router40;
	wire[`N2-1:0] out_router41;
	wire[`N2-1:0] out_router42;
	wire[`N2-1:0] out_router43;
	wire[`N2-1:0] out_router44;
	wire[`N2-1:0] out_router45;
	wire[`N2-1:0] out_router46;
	wire[`N2-1:0] out_router47;
	wire[`N2-1:0] out_router48;
	wire[`N2-1:0] out_router49;
	wire[`N2-1:0] out_router50;
	wire[`N2-1:0] out_router51;
	wire[`N2-1:0] out_router52;
	wire[`N2-1:0] out_router53;
	wire[`N2-1:0] out_router54;
	wire[`N2-1:0] out_router55;
	wire[`N2-1:0] out_router56;
	wire[`N2-1:0] out_router57;
	wire[`N2-1:0] out_router58;
	wire[`N2-1:0] out_router59;
	wire[`N2-1:0] out_router60;
	wire[`N2-1:0] out_router61;
	wire[`N2-1:0] out_router62;
	wire[`N2-1:0] out_router63;
	wire[`N2-1:0] out_router64;
	wire[`N2-1:0] out_router65;
	wire[`N2-1:0] out_router66;
	wire[`N2-1:0] out_router67;
	wire[`N2-1:0] out_router68;
	wire[`N2-1:0] out_router69;
	wire[`N2-1:0] out_router70;
	wire[`N2-1:0] out_router71;
	wire[`N2-1:0] out_router72;
	wire[`N2-1:0] out_router73;
	wire[`N2-1:0] out_router74;
	wire[`N2-1:0] out_router75;
	wire[`N2-1:0] out_router76;
	wire[`N2-1:0] out_router77;
	wire[`N2-1:0] out_router78;
	wire[`N2-1:0] out_router79;
	wire[`N2-1:0] out_router80;
	wire[`N2-1:0] out_router81;
	wire[`N2-1:0] out_router82;
	wire[`N2-1:0] out_router83;
	wire[`N2-1:0] out_router84;
	wire[`N2-1:0] out_router85;
	wire[`N2-1:0] out_router86;
	wire[`N2-1:0] out_router87;
	wire[`N2-1:0] out_router88;
	wire[`N2-1:0] out_router89;
	wire[`N2-1:0] out_router90;
	wire[`N2-1:0] out_router91;
	wire[`N2-1:0] out_router92;
	wire[`N2-1:0] out_router93;
	wire[`N2-1:0] out_router94;
	wire[`N2-1:0] out_router95;
	wire[`N2-1:0] out_router96;
	wire[`N2-1:0] out_router97;
	wire[`N2-1:0] out_router98;
	wire[`N2-1:0] out_router99;
	wire[`N2-1:0] out_router100;
	wire[`N2-1:0] out_router101;
	wire[`N2-1:0] out_router102;
	wire[`N2-1:0] out_router103;
	wire[`N2-1:0] out_router104;
	wire[`N2-1:0] out_router105;
	wire[`N2-1:0] out_router106;
	wire[`N2-1:0] out_router107;
	wire[`N2-1:0] out_router108;
	wire[`N2-1:0] out_router109;
	wire[`N2-1:0] out_router110;
	wire[`N2-1:0] out_router111;
	wire[`N2-1:0] out_router112;
	wire[`N2-1:0] out_router113;
	wire[`N2-1:0] out_router114;
	wire[`N2-1:0] out_router115;
	wire[`N2-1:0] out_router116;
	wire[`N2-1:0] out_router117;
	wire[`N2-1:0] out_router118;
	wire[`N2-1:0] out_router119;
	wire[`N2-1:0] out_router120;
	wire[`N2-1:0] out_router121;
	wire[`N2-1:0] out_router122;
	wire[`N2-1:0] out_router123;
	wire[`N2-1:0] out_router124;
	wire[`N2-1:0] out_router125;
	wire[`N2-1:0] out_router126;
	wire[`N2-1:0] out_router127;
	wire[`N2-1:0] out_router128;
	wire[`N2-1:0] out_router129;
	wire[`N2-1:0] out_router130;
	wire[`N2-1:0] out_router131;
	wire[`N2-1:0] out_router132;
	wire[`N2-1:0] out_router133;
	wire[`N2-1:0] out_router134;
	wire[`N2-1:0] out_router135;
	wire[`N2-1:0] out_router136;
	wire[`N2-1:0] out_router137;
	wire[`N2-1:0] out_router138;
	wire[`N2-1:0] out_router139;
	wire[`N2-1:0] out_router140;
	wire[`N2-1:0] out_router141;
	wire[`N2-1:0] out_router142;
	wire[`N2-1:0] out_router143;
	wire[`N2-1:0] out_router144;

	wire[`N2-1:0] r_min[0:`N_COUNT];	// в право по малой   образующей    данные от out_r1R
	wire[`N2-1:0] r_max[0:`N_COUNT];	// в право по большей образующей    данные от out_r2R
	wire[`N2-1:0] l_min[0:`N_COUNT];	// в лево  по малой   образующей    данные от out_r1L
	wire[`N2-1:0] l_max[0:`N_COUNT];	// в лево  по большей образующей    данные от out_r2L

	select_data_144 sel (.clk(clk), .sw_on(sw_on), .sw_sel_data(sw_sel_data), .sw_sel_router(sw_sel_router), .key_inc(key_inc), .key_dec(key_dec), .out_router1(out_router1), .out_router2(out_router2), .out_router3(out_router3), .out_router4(out_router4), .out_router5(out_router5), .out_router6(out_router6), .out_router7(out_router7), .out_router8(out_router8), .out_router9(out_router9), .out_router10(out_router10), .out_router11(out_router11), .out_router12(out_router12), .out_router13(out_router13), .out_router14(out_router14), .out_router15(out_router15), .out_router16(out_router16), .out_router17(out_router17), .out_router18(out_router18), .out_router19(out_router19), .out_router20(out_router20), .out_router21(out_router21), .out_router22(out_router22), .out_router23(out_router23), .out_router24(out_router24), .out_router25(out_router25), .out_router26(out_router26), .out_router27(out_router27), .out_router28(out_router28), .out_router29(out_router29), .out_router30(out_router30), .out_router31(out_router31), .out_router32(out_router32), .out_router33(out_router33), .out_router34(out_router34), .out_router35(out_router35), .out_router36(out_router36), .out_router37(out_router37), .out_router38(out_router38), .out_router39(out_router39), .out_router40(out_router40), .out_router41(out_router41), .out_router42(out_router42), .out_router43(out_router43), .out_router44(out_router44), .out_router45(out_router45), .out_router46(out_router46), .out_router47(out_router47), .out_router48(out_router48), .out_router49(out_router49), .out_router50(out_router50), .out_router51(out_router51), .out_router52(out_router52), .out_router53(out_router53), .out_router54(out_router54), .out_router55(out_router55), .out_router56(out_router56), .out_router57(out_router57), .out_router58(out_router58), .out_router59(out_router59), .out_router60(out_router60), .out_router61(out_router61), .out_router62(out_router62), .out_router63(out_router63), .out_router64(out_router64), .out_router65(out_router65), .out_router66(out_router66), .out_router67(out_router67), .out_router68(out_router68), .out_router69(out_router69), .out_router70(out_router70), .out_router71(out_router71), .out_router72(out_router72), .out_router73(out_router73), .out_router74(out_router74), .out_router75(out_router75), .out_router76(out_router76), .out_router77(out_router77), .out_router78(out_router78), .out_router79(out_router79), .out_router80(out_router80), .out_router81(out_router81), .out_router82(out_router82), .out_router83(out_router83), .out_router84(out_router84), .out_router85(out_router85), .out_router86(out_router86), .out_router87(out_router87), .out_router88(out_router88), .out_router89(out_router89), .out_router90(out_router90), .out_router91(out_router91), .out_router92(out_router92), .out_router93(out_router93), .out_router94(out_router94), .out_router95(out_router95), .out_router96(out_router96), .out_router97(out_router97), .out_router98(out_router98), .out_router99(out_router99), .out_router100(out_router100), .out_router101(out_router101), .out_router102(out_router102), .out_router103(out_router103), .out_router104(out_router104), .out_router105(out_router105), .out_router106(out_router106), .out_router107(out_router107), .out_router108(out_router108), .out_router109(out_router109), .out_router110(out_router110), .out_router111(out_router111), .out_router112(out_router112), .out_router113(out_router113), .out_router114(out_router114), .out_router115(out_router115), .out_router116(out_router116), .out_router117(out_router117), .out_router118(out_router118), .out_router119(out_router119), .out_router120(out_router120), .out_router121(out_router121), .out_router122(out_router122), .out_router123(out_router123), .out_router124(out_router124), .out_router125(out_router125), .out_router126(out_router126), .out_router127(out_router127), .out_router128(out_router128), .out_router129(out_router129), .out_router130(out_router130), .out_router131(out_router131), .out_router132(out_router132), .out_router133(out_router133), .out_router134(out_router134), .out_router135(out_router135), .out_router136(out_router136), .out_router137(out_router137), .out_router138(out_router138), .out_router139(out_router139), .out_router140(out_router140), .out_router141(out_router141), .out_router142(out_router142), .out_router143(out_router143), .out_router144(out_router144), .hex_data(hex_data), .hex_router(hex_router));

	apo_router_144_nodes r1 (.clk(clk), .router_name(8'b00000000), .in_free(out_router1), .in_r1R(l_min[8]), .in_r2R(l_max[9]), .in_r1L(r_min[136]), .in_r2L(r_max[135]), .out_r1R(r_min[0]), .out_r2R(r_max[0]), .out_r1L(l_min[0]), .out_r2L(l_max[0]), .out_data(out_data[0]));
	apo_router_144_nodes r2 (.clk(clk), .router_name(8'b00000001), .in_free(out_router2), .in_r1R(l_min[9]), .in_r2R(l_max[10]), .in_r1L(r_min[137]), .in_r2L(r_max[136]), .out_r1R(r_min[1]), .out_r2R(r_max[1]), .out_r1L(l_min[1]), .out_r2L(l_max[1]), .out_data(out_data[1]));
	apo_router_144_nodes r3 (.clk(clk), .router_name(8'b00000010), .in_free(out_router3), .in_r1R(l_min[10]), .in_r2R(l_max[11]), .in_r1L(r_min[138]), .in_r2L(r_max[137]), .out_r1R(r_min[2]), .out_r2R(r_max[2]), .out_r1L(l_min[2]), .out_r2L(l_max[2]), .out_data(out_data[2]));
	apo_router_144_nodes r4 (.clk(clk), .router_name(8'b00000011), .in_free(out_router4), .in_r1R(l_min[11]), .in_r2R(l_max[12]), .in_r1L(r_min[139]), .in_r2L(r_max[138]), .out_r1R(r_min[3]), .out_r2R(r_max[3]), .out_r1L(l_min[3]), .out_r2L(l_max[3]), .out_data(out_data[3]));
	apo_router_144_nodes r5 (.clk(clk), .router_name(8'b00000100), .in_free(out_router5), .in_r1R(l_min[12]), .in_r2R(l_max[13]), .in_r1L(r_min[140]), .in_r2L(r_max[139]), .out_r1R(r_min[4]), .out_r2R(r_max[4]), .out_r1L(l_min[4]), .out_r2L(l_max[4]), .out_data(out_data[4]));
	apo_router_144_nodes r6 (.clk(clk), .router_name(8'b00000101), .in_free(out_router6), .in_r1R(l_min[13]), .in_r2R(l_max[14]), .in_r1L(r_min[141]), .in_r2L(r_max[140]), .out_r1R(r_min[5]), .out_r2R(r_max[5]), .out_r1L(l_min[5]), .out_r2L(l_max[5]), .out_data(out_data[5]));
	apo_router_144_nodes r7 (.clk(clk), .router_name(8'b00000110), .in_free(out_router7), .in_r1R(l_min[14]), .in_r2R(l_max[15]), .in_r1L(r_min[142]), .in_r2L(r_max[141]), .out_r1R(r_min[6]), .out_r2R(r_max[6]), .out_r1L(l_min[6]), .out_r2L(l_max[6]), .out_data(out_data[6]));
	apo_router_144_nodes r8 (.clk(clk), .router_name(8'b00000111), .in_free(out_router8), .in_r1R(l_min[15]), .in_r2R(l_max[16]), .in_r1L(r_min[143]), .in_r2L(r_max[142]), .out_r1R(r_min[7]), .out_r2R(r_max[7]), .out_r1L(l_min[7]), .out_r2L(l_max[7]), .out_data(out_data[7]));
	apo_router_144_nodes r9 (.clk(clk), .router_name(8'b00001000), .in_free(out_router9), .in_r1R(l_min[16]), .in_r2R(l_max[17]), .in_r1L(r_min[0]), .in_r2L(r_max[143]), .out_r1R(r_min[8]), .out_r2R(r_max[8]), .out_r1L(l_min[8]), .out_r2L(l_max[8]), .out_data(out_data[8]));
	apo_router_144_nodes r10 (.clk(clk), .router_name(8'b00001001), .in_free(out_router10), .in_r1R(l_min[17]), .in_r2R(l_max[18]), .in_r1L(r_min[1]), .in_r2L(r_max[0]), .out_r1R(r_min[9]), .out_r2R(r_max[9]), .out_r1L(l_min[9]), .out_r2L(l_max[9]), .out_data(out_data[9]));
	apo_router_144_nodes r11 (.clk(clk), .router_name(8'b00001010), .in_free(out_router11), .in_r1R(l_min[18]), .in_r2R(l_max[19]), .in_r1L(r_min[2]), .in_r2L(r_max[1]), .out_r1R(r_min[10]), .out_r2R(r_max[10]), .out_r1L(l_min[10]), .out_r2L(l_max[10]), .out_data(out_data[10]));
	apo_router_144_nodes r12 (.clk(clk), .router_name(8'b00001011), .in_free(out_router12), .in_r1R(l_min[19]), .in_r2R(l_max[20]), .in_r1L(r_min[3]), .in_r2L(r_max[2]), .out_r1R(r_min[11]), .out_r2R(r_max[11]), .out_r1L(l_min[11]), .out_r2L(l_max[11]), .out_data(out_data[11]));
	apo_router_144_nodes r13 (.clk(clk), .router_name(8'b00001100), .in_free(out_router13), .in_r1R(l_min[20]), .in_r2R(l_max[21]), .in_r1L(r_min[4]), .in_r2L(r_max[3]), .out_r1R(r_min[12]), .out_r2R(r_max[12]), .out_r1L(l_min[12]), .out_r2L(l_max[12]), .out_data(out_data[12]));
	apo_router_144_nodes r14 (.clk(clk), .router_name(8'b00001101), .in_free(out_router14), .in_r1R(l_min[21]), .in_r2R(l_max[22]), .in_r1L(r_min[5]), .in_r2L(r_max[4]), .out_r1R(r_min[13]), .out_r2R(r_max[13]), .out_r1L(l_min[13]), .out_r2L(l_max[13]), .out_data(out_data[13]));
	apo_router_144_nodes r15 (.clk(clk), .router_name(8'b00001110), .in_free(out_router15), .in_r1R(l_min[22]), .in_r2R(l_max[23]), .in_r1L(r_min[6]), .in_r2L(r_max[5]), .out_r1R(r_min[14]), .out_r2R(r_max[14]), .out_r1L(l_min[14]), .out_r2L(l_max[14]), .out_data(out_data[14]));
	apo_router_144_nodes r16 (.clk(clk), .router_name(8'b00001111), .in_free(out_router16), .in_r1R(l_min[23]), .in_r2R(l_max[24]), .in_r1L(r_min[7]), .in_r2L(r_max[6]), .out_r1R(r_min[15]), .out_r2R(r_max[15]), .out_r1L(l_min[15]), .out_r2L(l_max[15]), .out_data(out_data[15]));
	apo_router_144_nodes r17 (.clk(clk), .router_name(8'b00010000), .in_free(out_router17), .in_r1R(l_min[24]), .in_r2R(l_max[25]), .in_r1L(r_min[8]), .in_r2L(r_max[7]), .out_r1R(r_min[16]), .out_r2R(r_max[16]), .out_r1L(l_min[16]), .out_r2L(l_max[16]), .out_data(out_data[16]));
	apo_router_144_nodes r18 (.clk(clk), .router_name(8'b00010001), .in_free(out_router18), .in_r1R(l_min[25]), .in_r2R(l_max[26]), .in_r1L(r_min[9]), .in_r2L(r_max[8]), .out_r1R(r_min[17]), .out_r2R(r_max[17]), .out_r1L(l_min[17]), .out_r2L(l_max[17]), .out_data(out_data[17]));
	apo_router_144_nodes r19 (.clk(clk), .router_name(8'b00010010), .in_free(out_router19), .in_r1R(l_min[26]), .in_r2R(l_max[27]), .in_r1L(r_min[10]), .in_r2L(r_max[9]), .out_r1R(r_min[18]), .out_r2R(r_max[18]), .out_r1L(l_min[18]), .out_r2L(l_max[18]), .out_data(out_data[18]));
	apo_router_144_nodes r20 (.clk(clk), .router_name(8'b00010011), .in_free(out_router20), .in_r1R(l_min[27]), .in_r2R(l_max[28]), .in_r1L(r_min[11]), .in_r2L(r_max[10]), .out_r1R(r_min[19]), .out_r2R(r_max[19]), .out_r1L(l_min[19]), .out_r2L(l_max[19]), .out_data(out_data[19]));
	apo_router_144_nodes r21 (.clk(clk), .router_name(8'b00010100), .in_free(out_router21), .in_r1R(l_min[28]), .in_r2R(l_max[29]), .in_r1L(r_min[12]), .in_r2L(r_max[11]), .out_r1R(r_min[20]), .out_r2R(r_max[20]), .out_r1L(l_min[20]), .out_r2L(l_max[20]), .out_data(out_data[20]));
	apo_router_144_nodes r22 (.clk(clk), .router_name(8'b00010101), .in_free(out_router22), .in_r1R(l_min[29]), .in_r2R(l_max[30]), .in_r1L(r_min[13]), .in_r2L(r_max[12]), .out_r1R(r_min[21]), .out_r2R(r_max[21]), .out_r1L(l_min[21]), .out_r2L(l_max[21]), .out_data(out_data[21]));
	apo_router_144_nodes r23 (.clk(clk), .router_name(8'b00010110), .in_free(out_router23), .in_r1R(l_min[30]), .in_r2R(l_max[31]), .in_r1L(r_min[14]), .in_r2L(r_max[13]), .out_r1R(r_min[22]), .out_r2R(r_max[22]), .out_r1L(l_min[22]), .out_r2L(l_max[22]), .out_data(out_data[22]));
	apo_router_144_nodes r24 (.clk(clk), .router_name(8'b00010111), .in_free(out_router24), .in_r1R(l_min[31]), .in_r2R(l_max[32]), .in_r1L(r_min[15]), .in_r2L(r_max[14]), .out_r1R(r_min[23]), .out_r2R(r_max[23]), .out_r1L(l_min[23]), .out_r2L(l_max[23]), .out_data(out_data[23]));
	apo_router_144_nodes r25 (.clk(clk), .router_name(8'b00011000), .in_free(out_router25), .in_r1R(l_min[32]), .in_r2R(l_max[33]), .in_r1L(r_min[16]), .in_r2L(r_max[15]), .out_r1R(r_min[24]), .out_r2R(r_max[24]), .out_r1L(l_min[24]), .out_r2L(l_max[24]), .out_data(out_data[24]));
	apo_router_144_nodes r26 (.clk(clk), .router_name(8'b00011001), .in_free(out_router26), .in_r1R(l_min[33]), .in_r2R(l_max[34]), .in_r1L(r_min[17]), .in_r2L(r_max[16]), .out_r1R(r_min[25]), .out_r2R(r_max[25]), .out_r1L(l_min[25]), .out_r2L(l_max[25]), .out_data(out_data[25]));
	apo_router_144_nodes r27 (.clk(clk), .router_name(8'b00011010), .in_free(out_router27), .in_r1R(l_min[34]), .in_r2R(l_max[35]), .in_r1L(r_min[18]), .in_r2L(r_max[17]), .out_r1R(r_min[26]), .out_r2R(r_max[26]), .out_r1L(l_min[26]), .out_r2L(l_max[26]), .out_data(out_data[26]));
	apo_router_144_nodes r28 (.clk(clk), .router_name(8'b00011011), .in_free(out_router28), .in_r1R(l_min[35]), .in_r2R(l_max[36]), .in_r1L(r_min[19]), .in_r2L(r_max[18]), .out_r1R(r_min[27]), .out_r2R(r_max[27]), .out_r1L(l_min[27]), .out_r2L(l_max[27]), .out_data(out_data[27]));
	apo_router_144_nodes r29 (.clk(clk), .router_name(8'b00011100), .in_free(out_router29), .in_r1R(l_min[36]), .in_r2R(l_max[37]), .in_r1L(r_min[20]), .in_r2L(r_max[19]), .out_r1R(r_min[28]), .out_r2R(r_max[28]), .out_r1L(l_min[28]), .out_r2L(l_max[28]), .out_data(out_data[28]));
	apo_router_144_nodes r30 (.clk(clk), .router_name(8'b00011101), .in_free(out_router30), .in_r1R(l_min[37]), .in_r2R(l_max[38]), .in_r1L(r_min[21]), .in_r2L(r_max[20]), .out_r1R(r_min[29]), .out_r2R(r_max[29]), .out_r1L(l_min[29]), .out_r2L(l_max[29]), .out_data(out_data[29]));
	apo_router_144_nodes r31 (.clk(clk), .router_name(8'b00011110), .in_free(out_router31), .in_r1R(l_min[38]), .in_r2R(l_max[39]), .in_r1L(r_min[22]), .in_r2L(r_max[21]), .out_r1R(r_min[30]), .out_r2R(r_max[30]), .out_r1L(l_min[30]), .out_r2L(l_max[30]), .out_data(out_data[30]));
	apo_router_144_nodes r32 (.clk(clk), .router_name(8'b00011111), .in_free(out_router32), .in_r1R(l_min[39]), .in_r2R(l_max[40]), .in_r1L(r_min[23]), .in_r2L(r_max[22]), .out_r1R(r_min[31]), .out_r2R(r_max[31]), .out_r1L(l_min[31]), .out_r2L(l_max[31]), .out_data(out_data[31]));
	apo_router_144_nodes r33 (.clk(clk), .router_name(8'b00100000), .in_free(out_router33), .in_r1R(l_min[40]), .in_r2R(l_max[41]), .in_r1L(r_min[24]), .in_r2L(r_max[23]), .out_r1R(r_min[32]), .out_r2R(r_max[32]), .out_r1L(l_min[32]), .out_r2L(l_max[32]), .out_data(out_data[32]));
	apo_router_144_nodes r34 (.clk(clk), .router_name(8'b00100001), .in_free(out_router34), .in_r1R(l_min[41]), .in_r2R(l_max[42]), .in_r1L(r_min[25]), .in_r2L(r_max[24]), .out_r1R(r_min[33]), .out_r2R(r_max[33]), .out_r1L(l_min[33]), .out_r2L(l_max[33]), .out_data(out_data[33]));
	apo_router_144_nodes r35 (.clk(clk), .router_name(8'b00100010), .in_free(out_router35), .in_r1R(l_min[42]), .in_r2R(l_max[43]), .in_r1L(r_min[26]), .in_r2L(r_max[25]), .out_r1R(r_min[34]), .out_r2R(r_max[34]), .out_r1L(l_min[34]), .out_r2L(l_max[34]), .out_data(out_data[34]));
	apo_router_144_nodes r36 (.clk(clk), .router_name(8'b00100011), .in_free(out_router36), .in_r1R(l_min[43]), .in_r2R(l_max[44]), .in_r1L(r_min[27]), .in_r2L(r_max[26]), .out_r1R(r_min[35]), .out_r2R(r_max[35]), .out_r1L(l_min[35]), .out_r2L(l_max[35]), .out_data(out_data[35]));
	apo_router_144_nodes r37 (.clk(clk), .router_name(8'b00100100), .in_free(out_router37), .in_r1R(l_min[44]), .in_r2R(l_max[45]), .in_r1L(r_min[28]), .in_r2L(r_max[27]), .out_r1R(r_min[36]), .out_r2R(r_max[36]), .out_r1L(l_min[36]), .out_r2L(l_max[36]), .out_data(out_data[36]));
	apo_router_144_nodes r38 (.clk(clk), .router_name(8'b00100101), .in_free(out_router38), .in_r1R(l_min[45]), .in_r2R(l_max[46]), .in_r1L(r_min[29]), .in_r2L(r_max[28]), .out_r1R(r_min[37]), .out_r2R(r_max[37]), .out_r1L(l_min[37]), .out_r2L(l_max[37]), .out_data(out_data[37]));
	apo_router_144_nodes r39 (.clk(clk), .router_name(8'b00100110), .in_free(out_router39), .in_r1R(l_min[46]), .in_r2R(l_max[47]), .in_r1L(r_min[30]), .in_r2L(r_max[29]), .out_r1R(r_min[38]), .out_r2R(r_max[38]), .out_r1L(l_min[38]), .out_r2L(l_max[38]), .out_data(out_data[38]));
	apo_router_144_nodes r40 (.clk(clk), .router_name(8'b00100111), .in_free(out_router40), .in_r1R(l_min[47]), .in_r2R(l_max[48]), .in_r1L(r_min[31]), .in_r2L(r_max[30]), .out_r1R(r_min[39]), .out_r2R(r_max[39]), .out_r1L(l_min[39]), .out_r2L(l_max[39]), .out_data(out_data[39]));
	apo_router_144_nodes r41 (.clk(clk), .router_name(8'b00101000), .in_free(out_router41), .in_r1R(l_min[48]), .in_r2R(l_max[49]), .in_r1L(r_min[32]), .in_r2L(r_max[31]), .out_r1R(r_min[40]), .out_r2R(r_max[40]), .out_r1L(l_min[40]), .out_r2L(l_max[40]), .out_data(out_data[40]));
	apo_router_144_nodes r42 (.clk(clk), .router_name(8'b00101001), .in_free(out_router42), .in_r1R(l_min[49]), .in_r2R(l_max[50]), .in_r1L(r_min[33]), .in_r2L(r_max[32]), .out_r1R(r_min[41]), .out_r2R(r_max[41]), .out_r1L(l_min[41]), .out_r2L(l_max[41]), .out_data(out_data[41]));
	apo_router_144_nodes r43 (.clk(clk), .router_name(8'b00101010), .in_free(out_router43), .in_r1R(l_min[50]), .in_r2R(l_max[51]), .in_r1L(r_min[34]), .in_r2L(r_max[33]), .out_r1R(r_min[42]), .out_r2R(r_max[42]), .out_r1L(l_min[42]), .out_r2L(l_max[42]), .out_data(out_data[42]));
	apo_router_144_nodes r44 (.clk(clk), .router_name(8'b00101011), .in_free(out_router44), .in_r1R(l_min[51]), .in_r2R(l_max[52]), .in_r1L(r_min[35]), .in_r2L(r_max[34]), .out_r1R(r_min[43]), .out_r2R(r_max[43]), .out_r1L(l_min[43]), .out_r2L(l_max[43]), .out_data(out_data[43]));
	apo_router_144_nodes r45 (.clk(clk), .router_name(8'b00101100), .in_free(out_router45), .in_r1R(l_min[52]), .in_r2R(l_max[53]), .in_r1L(r_min[36]), .in_r2L(r_max[35]), .out_r1R(r_min[44]), .out_r2R(r_max[44]), .out_r1L(l_min[44]), .out_r2L(l_max[44]), .out_data(out_data[44]));
	apo_router_144_nodes r46 (.clk(clk), .router_name(8'b00101101), .in_free(out_router46), .in_r1R(l_min[53]), .in_r2R(l_max[54]), .in_r1L(r_min[37]), .in_r2L(r_max[36]), .out_r1R(r_min[45]), .out_r2R(r_max[45]), .out_r1L(l_min[45]), .out_r2L(l_max[45]), .out_data(out_data[45]));
	apo_router_144_nodes r47 (.clk(clk), .router_name(8'b00101110), .in_free(out_router47), .in_r1R(l_min[54]), .in_r2R(l_max[55]), .in_r1L(r_min[38]), .in_r2L(r_max[37]), .out_r1R(r_min[46]), .out_r2R(r_max[46]), .out_r1L(l_min[46]), .out_r2L(l_max[46]), .out_data(out_data[46]));
	apo_router_144_nodes r48 (.clk(clk), .router_name(8'b00101111), .in_free(out_router48), .in_r1R(l_min[55]), .in_r2R(l_max[56]), .in_r1L(r_min[39]), .in_r2L(r_max[38]), .out_r1R(r_min[47]), .out_r2R(r_max[47]), .out_r1L(l_min[47]), .out_r2L(l_max[47]), .out_data(out_data[47]));
	apo_router_144_nodes r49 (.clk(clk), .router_name(8'b00110000), .in_free(out_router49), .in_r1R(l_min[56]), .in_r2R(l_max[57]), .in_r1L(r_min[40]), .in_r2L(r_max[39]), .out_r1R(r_min[48]), .out_r2R(r_max[48]), .out_r1L(l_min[48]), .out_r2L(l_max[48]), .out_data(out_data[48]));
	apo_router_144_nodes r50 (.clk(clk), .router_name(8'b00110001), .in_free(out_router50), .in_r1R(l_min[57]), .in_r2R(l_max[58]), .in_r1L(r_min[41]), .in_r2L(r_max[40]), .out_r1R(r_min[49]), .out_r2R(r_max[49]), .out_r1L(l_min[49]), .out_r2L(l_max[49]), .out_data(out_data[49]));
	apo_router_144_nodes r51 (.clk(clk), .router_name(8'b00110010), .in_free(out_router51), .in_r1R(l_min[58]), .in_r2R(l_max[59]), .in_r1L(r_min[42]), .in_r2L(r_max[41]), .out_r1R(r_min[50]), .out_r2R(r_max[50]), .out_r1L(l_min[50]), .out_r2L(l_max[50]), .out_data(out_data[50]));
	apo_router_144_nodes r52 (.clk(clk), .router_name(8'b00110011), .in_free(out_router52), .in_r1R(l_min[59]), .in_r2R(l_max[60]), .in_r1L(r_min[43]), .in_r2L(r_max[42]), .out_r1R(r_min[51]), .out_r2R(r_max[51]), .out_r1L(l_min[51]), .out_r2L(l_max[51]), .out_data(out_data[51]));
	apo_router_144_nodes r53 (.clk(clk), .router_name(8'b00110100), .in_free(out_router53), .in_r1R(l_min[60]), .in_r2R(l_max[61]), .in_r1L(r_min[44]), .in_r2L(r_max[43]), .out_r1R(r_min[52]), .out_r2R(r_max[52]), .out_r1L(l_min[52]), .out_r2L(l_max[52]), .out_data(out_data[52]));
	apo_router_144_nodes r54 (.clk(clk), .router_name(8'b00110101), .in_free(out_router54), .in_r1R(l_min[61]), .in_r2R(l_max[62]), .in_r1L(r_min[45]), .in_r2L(r_max[44]), .out_r1R(r_min[53]), .out_r2R(r_max[53]), .out_r1L(l_min[53]), .out_r2L(l_max[53]), .out_data(out_data[53]));
	apo_router_144_nodes r55 (.clk(clk), .router_name(8'b00110110), .in_free(out_router55), .in_r1R(l_min[62]), .in_r2R(l_max[63]), .in_r1L(r_min[46]), .in_r2L(r_max[45]), .out_r1R(r_min[54]), .out_r2R(r_max[54]), .out_r1L(l_min[54]), .out_r2L(l_max[54]), .out_data(out_data[54]));
	apo_router_144_nodes r56 (.clk(clk), .router_name(8'b00110111), .in_free(out_router56), .in_r1R(l_min[63]), .in_r2R(l_max[64]), .in_r1L(r_min[47]), .in_r2L(r_max[46]), .out_r1R(r_min[55]), .out_r2R(r_max[55]), .out_r1L(l_min[55]), .out_r2L(l_max[55]), .out_data(out_data[55]));
	apo_router_144_nodes r57 (.clk(clk), .router_name(8'b00111000), .in_free(out_router57), .in_r1R(l_min[64]), .in_r2R(l_max[65]), .in_r1L(r_min[48]), .in_r2L(r_max[47]), .out_r1R(r_min[56]), .out_r2R(r_max[56]), .out_r1L(l_min[56]), .out_r2L(l_max[56]), .out_data(out_data[56]));
	apo_router_144_nodes r58 (.clk(clk), .router_name(8'b00111001), .in_free(out_router58), .in_r1R(l_min[65]), .in_r2R(l_max[66]), .in_r1L(r_min[49]), .in_r2L(r_max[48]), .out_r1R(r_min[57]), .out_r2R(r_max[57]), .out_r1L(l_min[57]), .out_r2L(l_max[57]), .out_data(out_data[57]));
	apo_router_144_nodes r59 (.clk(clk), .router_name(8'b00111010), .in_free(out_router59), .in_r1R(l_min[66]), .in_r2R(l_max[67]), .in_r1L(r_min[50]), .in_r2L(r_max[49]), .out_r1R(r_min[58]), .out_r2R(r_max[58]), .out_r1L(l_min[58]), .out_r2L(l_max[58]), .out_data(out_data[58]));
	apo_router_144_nodes r60 (.clk(clk), .router_name(8'b00111011), .in_free(out_router60), .in_r1R(l_min[67]), .in_r2R(l_max[68]), .in_r1L(r_min[51]), .in_r2L(r_max[50]), .out_r1R(r_min[59]), .out_r2R(r_max[59]), .out_r1L(l_min[59]), .out_r2L(l_max[59]), .out_data(out_data[59]));
	apo_router_144_nodes r61 (.clk(clk), .router_name(8'b00111100), .in_free(out_router61), .in_r1R(l_min[68]), .in_r2R(l_max[69]), .in_r1L(r_min[52]), .in_r2L(r_max[51]), .out_r1R(r_min[60]), .out_r2R(r_max[60]), .out_r1L(l_min[60]), .out_r2L(l_max[60]), .out_data(out_data[60]));
	apo_router_144_nodes r62 (.clk(clk), .router_name(8'b00111101), .in_free(out_router62), .in_r1R(l_min[69]), .in_r2R(l_max[70]), .in_r1L(r_min[53]), .in_r2L(r_max[52]), .out_r1R(r_min[61]), .out_r2R(r_max[61]), .out_r1L(l_min[61]), .out_r2L(l_max[61]), .out_data(out_data[61]));
	apo_router_144_nodes r63 (.clk(clk), .router_name(8'b00111110), .in_free(out_router63), .in_r1R(l_min[70]), .in_r2R(l_max[71]), .in_r1L(r_min[54]), .in_r2L(r_max[53]), .out_r1R(r_min[62]), .out_r2R(r_max[62]), .out_r1L(l_min[62]), .out_r2L(l_max[62]), .out_data(out_data[62]));
	apo_router_144_nodes r64 (.clk(clk), .router_name(8'b00111111), .in_free(out_router64), .in_r1R(l_min[71]), .in_r2R(l_max[72]), .in_r1L(r_min[55]), .in_r2L(r_max[54]), .out_r1R(r_min[63]), .out_r2R(r_max[63]), .out_r1L(l_min[63]), .out_r2L(l_max[63]), .out_data(out_data[63]));
	apo_router_144_nodes r65 (.clk(clk), .router_name(8'b01000000), .in_free(out_router65), .in_r1R(l_min[72]), .in_r2R(l_max[73]), .in_r1L(r_min[56]), .in_r2L(r_max[55]), .out_r1R(r_min[64]), .out_r2R(r_max[64]), .out_r1L(l_min[64]), .out_r2L(l_max[64]), .out_data(out_data[64]));
	apo_router_144_nodes r66 (.clk(clk), .router_name(8'b01000001), .in_free(out_router66), .in_r1R(l_min[73]), .in_r2R(l_max[74]), .in_r1L(r_min[57]), .in_r2L(r_max[56]), .out_r1R(r_min[65]), .out_r2R(r_max[65]), .out_r1L(l_min[65]), .out_r2L(l_max[65]), .out_data(out_data[65]));
	apo_router_144_nodes r67 (.clk(clk), .router_name(8'b01000010), .in_free(out_router67), .in_r1R(l_min[74]), .in_r2R(l_max[75]), .in_r1L(r_min[58]), .in_r2L(r_max[57]), .out_r1R(r_min[66]), .out_r2R(r_max[66]), .out_r1L(l_min[66]), .out_r2L(l_max[66]), .out_data(out_data[66]));
	apo_router_144_nodes r68 (.clk(clk), .router_name(8'b01000011), .in_free(out_router68), .in_r1R(l_min[75]), .in_r2R(l_max[76]), .in_r1L(r_min[59]), .in_r2L(r_max[58]), .out_r1R(r_min[67]), .out_r2R(r_max[67]), .out_r1L(l_min[67]), .out_r2L(l_max[67]), .out_data(out_data[67]));
	apo_router_144_nodes r69 (.clk(clk), .router_name(8'b01000100), .in_free(out_router69), .in_r1R(l_min[76]), .in_r2R(l_max[77]), .in_r1L(r_min[60]), .in_r2L(r_max[59]), .out_r1R(r_min[68]), .out_r2R(r_max[68]), .out_r1L(l_min[68]), .out_r2L(l_max[68]), .out_data(out_data[68]));
	apo_router_144_nodes r70 (.clk(clk), .router_name(8'b01000101), .in_free(out_router70), .in_r1R(l_min[77]), .in_r2R(l_max[78]), .in_r1L(r_min[61]), .in_r2L(r_max[60]), .out_r1R(r_min[69]), .out_r2R(r_max[69]), .out_r1L(l_min[69]), .out_r2L(l_max[69]), .out_data(out_data[69]));
	apo_router_144_nodes r71 (.clk(clk), .router_name(8'b01000110), .in_free(out_router71), .in_r1R(l_min[78]), .in_r2R(l_max[79]), .in_r1L(r_min[62]), .in_r2L(r_max[61]), .out_r1R(r_min[70]), .out_r2R(r_max[70]), .out_r1L(l_min[70]), .out_r2L(l_max[70]), .out_data(out_data[70]));
	apo_router_144_nodes r72 (.clk(clk), .router_name(8'b01000111), .in_free(out_router72), .in_r1R(l_min[79]), .in_r2R(l_max[80]), .in_r1L(r_min[63]), .in_r2L(r_max[62]), .out_r1R(r_min[71]), .out_r2R(r_max[71]), .out_r1L(l_min[71]), .out_r2L(l_max[71]), .out_data(out_data[71]));
	apo_router_144_nodes r73 (.clk(clk), .router_name(8'b01001000), .in_free(out_router73), .in_r1R(l_min[80]), .in_r2R(l_max[81]), .in_r1L(r_min[64]), .in_r2L(r_max[63]), .out_r1R(r_min[72]), .out_r2R(r_max[72]), .out_r1L(l_min[72]), .out_r2L(l_max[72]), .out_data(out_data[72]));
	apo_router_144_nodes r74 (.clk(clk), .router_name(8'b01001001), .in_free(out_router74), .in_r1R(l_min[81]), .in_r2R(l_max[82]), .in_r1L(r_min[65]), .in_r2L(r_max[64]), .out_r1R(r_min[73]), .out_r2R(r_max[73]), .out_r1L(l_min[73]), .out_r2L(l_max[73]), .out_data(out_data[73]));
	apo_router_144_nodes r75 (.clk(clk), .router_name(8'b01001010), .in_free(out_router75), .in_r1R(l_min[82]), .in_r2R(l_max[83]), .in_r1L(r_min[66]), .in_r2L(r_max[65]), .out_r1R(r_min[74]), .out_r2R(r_max[74]), .out_r1L(l_min[74]), .out_r2L(l_max[74]), .out_data(out_data[74]));
	apo_router_144_nodes r76 (.clk(clk), .router_name(8'b01001011), .in_free(out_router76), .in_r1R(l_min[83]), .in_r2R(l_max[84]), .in_r1L(r_min[67]), .in_r2L(r_max[66]), .out_r1R(r_min[75]), .out_r2R(r_max[75]), .out_r1L(l_min[75]), .out_r2L(l_max[75]), .out_data(out_data[75]));
	apo_router_144_nodes r77 (.clk(clk), .router_name(8'b01001100), .in_free(out_router77), .in_r1R(l_min[84]), .in_r2R(l_max[85]), .in_r1L(r_min[68]), .in_r2L(r_max[67]), .out_r1R(r_min[76]), .out_r2R(r_max[76]), .out_r1L(l_min[76]), .out_r2L(l_max[76]), .out_data(out_data[76]));
	apo_router_144_nodes r78 (.clk(clk), .router_name(8'b01001101), .in_free(out_router78), .in_r1R(l_min[85]), .in_r2R(l_max[86]), .in_r1L(r_min[69]), .in_r2L(r_max[68]), .out_r1R(r_min[77]), .out_r2R(r_max[77]), .out_r1L(l_min[77]), .out_r2L(l_max[77]), .out_data(out_data[77]));
	apo_router_144_nodes r79 (.clk(clk), .router_name(8'b01001110), .in_free(out_router79), .in_r1R(l_min[86]), .in_r2R(l_max[87]), .in_r1L(r_min[70]), .in_r2L(r_max[69]), .out_r1R(r_min[78]), .out_r2R(r_max[78]), .out_r1L(l_min[78]), .out_r2L(l_max[78]), .out_data(out_data[78]));
	apo_router_144_nodes r80 (.clk(clk), .router_name(8'b01001111), .in_free(out_router80), .in_r1R(l_min[87]), .in_r2R(l_max[88]), .in_r1L(r_min[71]), .in_r2L(r_max[70]), .out_r1R(r_min[79]), .out_r2R(r_max[79]), .out_r1L(l_min[79]), .out_r2L(l_max[79]), .out_data(out_data[79]));
	apo_router_144_nodes r81 (.clk(clk), .router_name(8'b01010000), .in_free(out_router81), .in_r1R(l_min[88]), .in_r2R(l_max[89]), .in_r1L(r_min[72]), .in_r2L(r_max[71]), .out_r1R(r_min[80]), .out_r2R(r_max[80]), .out_r1L(l_min[80]), .out_r2L(l_max[80]), .out_data(out_data[80]));
	apo_router_144_nodes r82 (.clk(clk), .router_name(8'b01010001), .in_free(out_router82), .in_r1R(l_min[89]), .in_r2R(l_max[90]), .in_r1L(r_min[73]), .in_r2L(r_max[72]), .out_r1R(r_min[81]), .out_r2R(r_max[81]), .out_r1L(l_min[81]), .out_r2L(l_max[81]), .out_data(out_data[81]));
	apo_router_144_nodes r83 (.clk(clk), .router_name(8'b01010010), .in_free(out_router83), .in_r1R(l_min[90]), .in_r2R(l_max[91]), .in_r1L(r_min[74]), .in_r2L(r_max[73]), .out_r1R(r_min[82]), .out_r2R(r_max[82]), .out_r1L(l_min[82]), .out_r2L(l_max[82]), .out_data(out_data[82]));
	apo_router_144_nodes r84 (.clk(clk), .router_name(8'b01010011), .in_free(out_router84), .in_r1R(l_min[91]), .in_r2R(l_max[92]), .in_r1L(r_min[75]), .in_r2L(r_max[74]), .out_r1R(r_min[83]), .out_r2R(r_max[83]), .out_r1L(l_min[83]), .out_r2L(l_max[83]), .out_data(out_data[83]));
	apo_router_144_nodes r85 (.clk(clk), .router_name(8'b01010100), .in_free(out_router85), .in_r1R(l_min[92]), .in_r2R(l_max[93]), .in_r1L(r_min[76]), .in_r2L(r_max[75]), .out_r1R(r_min[84]), .out_r2R(r_max[84]), .out_r1L(l_min[84]), .out_r2L(l_max[84]), .out_data(out_data[84]));
	apo_router_144_nodes r86 (.clk(clk), .router_name(8'b01010101), .in_free(out_router86), .in_r1R(l_min[93]), .in_r2R(l_max[94]), .in_r1L(r_min[77]), .in_r2L(r_max[76]), .out_r1R(r_min[85]), .out_r2R(r_max[85]), .out_r1L(l_min[85]), .out_r2L(l_max[85]), .out_data(out_data[85]));
	apo_router_144_nodes r87 (.clk(clk), .router_name(8'b01010110), .in_free(out_router87), .in_r1R(l_min[94]), .in_r2R(l_max[95]), .in_r1L(r_min[78]), .in_r2L(r_max[77]), .out_r1R(r_min[86]), .out_r2R(r_max[86]), .out_r1L(l_min[86]), .out_r2L(l_max[86]), .out_data(out_data[86]));
	apo_router_144_nodes r88 (.clk(clk), .router_name(8'b01010111), .in_free(out_router88), .in_r1R(l_min[95]), .in_r2R(l_max[96]), .in_r1L(r_min[79]), .in_r2L(r_max[78]), .out_r1R(r_min[87]), .out_r2R(r_max[87]), .out_r1L(l_min[87]), .out_r2L(l_max[87]), .out_data(out_data[87]));
	apo_router_144_nodes r89 (.clk(clk), .router_name(8'b01011000), .in_free(out_router89), .in_r1R(l_min[96]), .in_r2R(l_max[97]), .in_r1L(r_min[80]), .in_r2L(r_max[79]), .out_r1R(r_min[88]), .out_r2R(r_max[88]), .out_r1L(l_min[88]), .out_r2L(l_max[88]), .out_data(out_data[88]));
	apo_router_144_nodes r90 (.clk(clk), .router_name(8'b01011001), .in_free(out_router90), .in_r1R(l_min[97]), .in_r2R(l_max[98]), .in_r1L(r_min[81]), .in_r2L(r_max[80]), .out_r1R(r_min[89]), .out_r2R(r_max[89]), .out_r1L(l_min[89]), .out_r2L(l_max[89]), .out_data(out_data[89]));
	apo_router_144_nodes r91 (.clk(clk), .router_name(8'b01011010), .in_free(out_router91), .in_r1R(l_min[98]), .in_r2R(l_max[99]), .in_r1L(r_min[82]), .in_r2L(r_max[81]), .out_r1R(r_min[90]), .out_r2R(r_max[90]), .out_r1L(l_min[90]), .out_r2L(l_max[90]), .out_data(out_data[90]));
	apo_router_144_nodes r92 (.clk(clk), .router_name(8'b01011011), .in_free(out_router92), .in_r1R(l_min[99]), .in_r2R(l_max[100]), .in_r1L(r_min[83]), .in_r2L(r_max[82]), .out_r1R(r_min[91]), .out_r2R(r_max[91]), .out_r1L(l_min[91]), .out_r2L(l_max[91]), .out_data(out_data[91]));
	apo_router_144_nodes r93 (.clk(clk), .router_name(8'b01011100), .in_free(out_router93), .in_r1R(l_min[100]), .in_r2R(l_max[101]), .in_r1L(r_min[84]), .in_r2L(r_max[83]), .out_r1R(r_min[92]), .out_r2R(r_max[92]), .out_r1L(l_min[92]), .out_r2L(l_max[92]), .out_data(out_data[92]));
	apo_router_144_nodes r94 (.clk(clk), .router_name(8'b01011101), .in_free(out_router94), .in_r1R(l_min[101]), .in_r2R(l_max[102]), .in_r1L(r_min[85]), .in_r2L(r_max[84]), .out_r1R(r_min[93]), .out_r2R(r_max[93]), .out_r1L(l_min[93]), .out_r2L(l_max[93]), .out_data(out_data[93]));
	apo_router_144_nodes r95 (.clk(clk), .router_name(8'b01011110), .in_free(out_router95), .in_r1R(l_min[102]), .in_r2R(l_max[103]), .in_r1L(r_min[86]), .in_r2L(r_max[85]), .out_r1R(r_min[94]), .out_r2R(r_max[94]), .out_r1L(l_min[94]), .out_r2L(l_max[94]), .out_data(out_data[94]));
	apo_router_144_nodes r96 (.clk(clk), .router_name(8'b01011111), .in_free(out_router96), .in_r1R(l_min[103]), .in_r2R(l_max[104]), .in_r1L(r_min[87]), .in_r2L(r_max[86]), .out_r1R(r_min[95]), .out_r2R(r_max[95]), .out_r1L(l_min[95]), .out_r2L(l_max[95]), .out_data(out_data[95]));
	apo_router_144_nodes r97 (.clk(clk), .router_name(8'b01100000), .in_free(out_router97), .in_r1R(l_min[104]), .in_r2R(l_max[105]), .in_r1L(r_min[88]), .in_r2L(r_max[87]), .out_r1R(r_min[96]), .out_r2R(r_max[96]), .out_r1L(l_min[96]), .out_r2L(l_max[96]), .out_data(out_data[96]));
	apo_router_144_nodes r98 (.clk(clk), .router_name(8'b01100001), .in_free(out_router98), .in_r1R(l_min[105]), .in_r2R(l_max[106]), .in_r1L(r_min[89]), .in_r2L(r_max[88]), .out_r1R(r_min[97]), .out_r2R(r_max[97]), .out_r1L(l_min[97]), .out_r2L(l_max[97]), .out_data(out_data[97]));
	apo_router_144_nodes r99 (.clk(clk), .router_name(8'b01100010), .in_free(out_router99), .in_r1R(l_min[106]), .in_r2R(l_max[107]), .in_r1L(r_min[90]), .in_r2L(r_max[89]), .out_r1R(r_min[98]), .out_r2R(r_max[98]), .out_r1L(l_min[98]), .out_r2L(l_max[98]), .out_data(out_data[98]));
	apo_router_144_nodes r100 (.clk(clk), .router_name(8'b01100011), .in_free(out_router100), .in_r1R(l_min[107]), .in_r2R(l_max[108]), .in_r1L(r_min[91]), .in_r2L(r_max[90]), .out_r1R(r_min[99]), .out_r2R(r_max[99]), .out_r1L(l_min[99]), .out_r2L(l_max[99]), .out_data(out_data[99]));
	apo_router_144_nodes r101 (.clk(clk), .router_name(8'b01100100), .in_free(out_router101), .in_r1R(l_min[108]), .in_r2R(l_max[109]), .in_r1L(r_min[92]), .in_r2L(r_max[91]), .out_r1R(r_min[100]), .out_r2R(r_max[100]), .out_r1L(l_min[100]), .out_r2L(l_max[100]), .out_data(out_data[100]));
	apo_router_144_nodes r102 (.clk(clk), .router_name(8'b01100101), .in_free(out_router102), .in_r1R(l_min[109]), .in_r2R(l_max[110]), .in_r1L(r_min[93]), .in_r2L(r_max[92]), .out_r1R(r_min[101]), .out_r2R(r_max[101]), .out_r1L(l_min[101]), .out_r2L(l_max[101]), .out_data(out_data[101]));
	apo_router_144_nodes r103 (.clk(clk), .router_name(8'b01100110), .in_free(out_router103), .in_r1R(l_min[110]), .in_r2R(l_max[111]), .in_r1L(r_min[94]), .in_r2L(r_max[93]), .out_r1R(r_min[102]), .out_r2R(r_max[102]), .out_r1L(l_min[102]), .out_r2L(l_max[102]), .out_data(out_data[102]));
	apo_router_144_nodes r104 (.clk(clk), .router_name(8'b01100111), .in_free(out_router104), .in_r1R(l_min[111]), .in_r2R(l_max[112]), .in_r1L(r_min[95]), .in_r2L(r_max[94]), .out_r1R(r_min[103]), .out_r2R(r_max[103]), .out_r1L(l_min[103]), .out_r2L(l_max[103]), .out_data(out_data[103]));
	apo_router_144_nodes r105 (.clk(clk), .router_name(8'b01101000), .in_free(out_router105), .in_r1R(l_min[112]), .in_r2R(l_max[113]), .in_r1L(r_min[96]), .in_r2L(r_max[95]), .out_r1R(r_min[104]), .out_r2R(r_max[104]), .out_r1L(l_min[104]), .out_r2L(l_max[104]), .out_data(out_data[104]));
	apo_router_144_nodes r106 (.clk(clk), .router_name(8'b01101001), .in_free(out_router106), .in_r1R(l_min[113]), .in_r2R(l_max[114]), .in_r1L(r_min[97]), .in_r2L(r_max[96]), .out_r1R(r_min[105]), .out_r2R(r_max[105]), .out_r1L(l_min[105]), .out_r2L(l_max[105]), .out_data(out_data[105]));
	apo_router_144_nodes r107 (.clk(clk), .router_name(8'b01101010), .in_free(out_router107), .in_r1R(l_min[114]), .in_r2R(l_max[115]), .in_r1L(r_min[98]), .in_r2L(r_max[97]), .out_r1R(r_min[106]), .out_r2R(r_max[106]), .out_r1L(l_min[106]), .out_r2L(l_max[106]), .out_data(out_data[106]));
	apo_router_144_nodes r108 (.clk(clk), .router_name(8'b01101011), .in_free(out_router108), .in_r1R(l_min[115]), .in_r2R(l_max[116]), .in_r1L(r_min[99]), .in_r2L(r_max[98]), .out_r1R(r_min[107]), .out_r2R(r_max[107]), .out_r1L(l_min[107]), .out_r2L(l_max[107]), .out_data(out_data[107]));
	apo_router_144_nodes r109 (.clk(clk), .router_name(8'b01101100), .in_free(out_router109), .in_r1R(l_min[116]), .in_r2R(l_max[117]), .in_r1L(r_min[100]), .in_r2L(r_max[99]), .out_r1R(r_min[108]), .out_r2R(r_max[108]), .out_r1L(l_min[108]), .out_r2L(l_max[108]), .out_data(out_data[108]));
	apo_router_144_nodes r110 (.clk(clk), .router_name(8'b01101101), .in_free(out_router110), .in_r1R(l_min[117]), .in_r2R(l_max[118]), .in_r1L(r_min[101]), .in_r2L(r_max[100]), .out_r1R(r_min[109]), .out_r2R(r_max[109]), .out_r1L(l_min[109]), .out_r2L(l_max[109]), .out_data(out_data[109]));
	apo_router_144_nodes r111 (.clk(clk), .router_name(8'b01101110), .in_free(out_router111), .in_r1R(l_min[118]), .in_r2R(l_max[119]), .in_r1L(r_min[102]), .in_r2L(r_max[101]), .out_r1R(r_min[110]), .out_r2R(r_max[110]), .out_r1L(l_min[110]), .out_r2L(l_max[110]), .out_data(out_data[110]));
	apo_router_144_nodes r112 (.clk(clk), .router_name(8'b01101111), .in_free(out_router112), .in_r1R(l_min[119]), .in_r2R(l_max[120]), .in_r1L(r_min[103]), .in_r2L(r_max[102]), .out_r1R(r_min[111]), .out_r2R(r_max[111]), .out_r1L(l_min[111]), .out_r2L(l_max[111]), .out_data(out_data[111]));
	apo_router_144_nodes r113 (.clk(clk), .router_name(8'b01110000), .in_free(out_router113), .in_r1R(l_min[120]), .in_r2R(l_max[121]), .in_r1L(r_min[104]), .in_r2L(r_max[103]), .out_r1R(r_min[112]), .out_r2R(r_max[112]), .out_r1L(l_min[112]), .out_r2L(l_max[112]), .out_data(out_data[112]));
	apo_router_144_nodes r114 (.clk(clk), .router_name(8'b01110001), .in_free(out_router114), .in_r1R(l_min[121]), .in_r2R(l_max[122]), .in_r1L(r_min[105]), .in_r2L(r_max[104]), .out_r1R(r_min[113]), .out_r2R(r_max[113]), .out_r1L(l_min[113]), .out_r2L(l_max[113]), .out_data(out_data[113]));
	apo_router_144_nodes r115 (.clk(clk), .router_name(8'b01110010), .in_free(out_router115), .in_r1R(l_min[122]), .in_r2R(l_max[123]), .in_r1L(r_min[106]), .in_r2L(r_max[105]), .out_r1R(r_min[114]), .out_r2R(r_max[114]), .out_r1L(l_min[114]), .out_r2L(l_max[114]), .out_data(out_data[114]));
	apo_router_144_nodes r116 (.clk(clk), .router_name(8'b01110011), .in_free(out_router116), .in_r1R(l_min[123]), .in_r2R(l_max[124]), .in_r1L(r_min[107]), .in_r2L(r_max[106]), .out_r1R(r_min[115]), .out_r2R(r_max[115]), .out_r1L(l_min[115]), .out_r2L(l_max[115]), .out_data(out_data[115]));
	apo_router_144_nodes r117 (.clk(clk), .router_name(8'b01110100), .in_free(out_router117), .in_r1R(l_min[124]), .in_r2R(l_max[125]), .in_r1L(r_min[108]), .in_r2L(r_max[107]), .out_r1R(r_min[116]), .out_r2R(r_max[116]), .out_r1L(l_min[116]), .out_r2L(l_max[116]), .out_data(out_data[116]));
	apo_router_144_nodes r118 (.clk(clk), .router_name(8'b01110101), .in_free(out_router118), .in_r1R(l_min[125]), .in_r2R(l_max[126]), .in_r1L(r_min[109]), .in_r2L(r_max[108]), .out_r1R(r_min[117]), .out_r2R(r_max[117]), .out_r1L(l_min[117]), .out_r2L(l_max[117]), .out_data(out_data[117]));
	apo_router_144_nodes r119 (.clk(clk), .router_name(8'b01110110), .in_free(out_router119), .in_r1R(l_min[126]), .in_r2R(l_max[127]), .in_r1L(r_min[110]), .in_r2L(r_max[109]), .out_r1R(r_min[118]), .out_r2R(r_max[118]), .out_r1L(l_min[118]), .out_r2L(l_max[118]), .out_data(out_data[118]));
	apo_router_144_nodes r120 (.clk(clk), .router_name(8'b01110111), .in_free(out_router120), .in_r1R(l_min[127]), .in_r2R(l_max[128]), .in_r1L(r_min[111]), .in_r2L(r_max[110]), .out_r1R(r_min[119]), .out_r2R(r_max[119]), .out_r1L(l_min[119]), .out_r2L(l_max[119]), .out_data(out_data[119]));
	apo_router_144_nodes r121 (.clk(clk), .router_name(8'b01111000), .in_free(out_router121), .in_r1R(l_min[128]), .in_r2R(l_max[129]), .in_r1L(r_min[112]), .in_r2L(r_max[111]), .out_r1R(r_min[120]), .out_r2R(r_max[120]), .out_r1L(l_min[120]), .out_r2L(l_max[120]), .out_data(out_data[120]));
	apo_router_144_nodes r122 (.clk(clk), .router_name(8'b01111001), .in_free(out_router122), .in_r1R(l_min[129]), .in_r2R(l_max[130]), .in_r1L(r_min[113]), .in_r2L(r_max[112]), .out_r1R(r_min[121]), .out_r2R(r_max[121]), .out_r1L(l_min[121]), .out_r2L(l_max[121]), .out_data(out_data[121]));
	apo_router_144_nodes r123 (.clk(clk), .router_name(8'b01111010), .in_free(out_router123), .in_r1R(l_min[130]), .in_r2R(l_max[131]), .in_r1L(r_min[114]), .in_r2L(r_max[113]), .out_r1R(r_min[122]), .out_r2R(r_max[122]), .out_r1L(l_min[122]), .out_r2L(l_max[122]), .out_data(out_data[122]));
	apo_router_144_nodes r124 (.clk(clk), .router_name(8'b01111011), .in_free(out_router124), .in_r1R(l_min[131]), .in_r2R(l_max[132]), .in_r1L(r_min[115]), .in_r2L(r_max[114]), .out_r1R(r_min[123]), .out_r2R(r_max[123]), .out_r1L(l_min[123]), .out_r2L(l_max[123]), .out_data(out_data[123]));
	apo_router_144_nodes r125 (.clk(clk), .router_name(8'b01111100), .in_free(out_router125), .in_r1R(l_min[132]), .in_r2R(l_max[133]), .in_r1L(r_min[116]), .in_r2L(r_max[115]), .out_r1R(r_min[124]), .out_r2R(r_max[124]), .out_r1L(l_min[124]), .out_r2L(l_max[124]), .out_data(out_data[124]));
	apo_router_144_nodes r126 (.clk(clk), .router_name(8'b01111101), .in_free(out_router126), .in_r1R(l_min[133]), .in_r2R(l_max[134]), .in_r1L(r_min[117]), .in_r2L(r_max[116]), .out_r1R(r_min[125]), .out_r2R(r_max[125]), .out_r1L(l_min[125]), .out_r2L(l_max[125]), .out_data(out_data[125]));
	apo_router_144_nodes r127 (.clk(clk), .router_name(8'b01111110), .in_free(out_router127), .in_r1R(l_min[134]), .in_r2R(l_max[135]), .in_r1L(r_min[118]), .in_r2L(r_max[117]), .out_r1R(r_min[126]), .out_r2R(r_max[126]), .out_r1L(l_min[126]), .out_r2L(l_max[126]), .out_data(out_data[126]));
	apo_router_144_nodes r128 (.clk(clk), .router_name(8'b01111111), .in_free(out_router128), .in_r1R(l_min[135]), .in_r2R(l_max[136]), .in_r1L(r_min[119]), .in_r2L(r_max[118]), .out_r1R(r_min[127]), .out_r2R(r_max[127]), .out_r1L(l_min[127]), .out_r2L(l_max[127]), .out_data(out_data[127]));
	apo_router_144_nodes r129 (.clk(clk), .router_name(8'b10000000), .in_free(out_router129), .in_r1R(l_min[136]), .in_r2R(l_max[137]), .in_r1L(r_min[120]), .in_r2L(r_max[119]), .out_r1R(r_min[128]), .out_r2R(r_max[128]), .out_r1L(l_min[128]), .out_r2L(l_max[128]), .out_data(out_data[128]));
	apo_router_144_nodes r130 (.clk(clk), .router_name(8'b10000001), .in_free(out_router130), .in_r1R(l_min[137]), .in_r2R(l_max[138]), .in_r1L(r_min[121]), .in_r2L(r_max[120]), .out_r1R(r_min[129]), .out_r2R(r_max[129]), .out_r1L(l_min[129]), .out_r2L(l_max[129]), .out_data(out_data[129]));
	apo_router_144_nodes r131 (.clk(clk), .router_name(8'b10000010), .in_free(out_router131), .in_r1R(l_min[138]), .in_r2R(l_max[139]), .in_r1L(r_min[122]), .in_r2L(r_max[121]), .out_r1R(r_min[130]), .out_r2R(r_max[130]), .out_r1L(l_min[130]), .out_r2L(l_max[130]), .out_data(out_data[130]));
	apo_router_144_nodes r132 (.clk(clk), .router_name(8'b10000011), .in_free(out_router132), .in_r1R(l_min[139]), .in_r2R(l_max[140]), .in_r1L(r_min[123]), .in_r2L(r_max[122]), .out_r1R(r_min[131]), .out_r2R(r_max[131]), .out_r1L(l_min[131]), .out_r2L(l_max[131]), .out_data(out_data[131]));
	apo_router_144_nodes r133 (.clk(clk), .router_name(8'b10000100), .in_free(out_router133), .in_r1R(l_min[140]), .in_r2R(l_max[141]), .in_r1L(r_min[124]), .in_r2L(r_max[123]), .out_r1R(r_min[132]), .out_r2R(r_max[132]), .out_r1L(l_min[132]), .out_r2L(l_max[132]), .out_data(out_data[132]));
	apo_router_144_nodes r134 (.clk(clk), .router_name(8'b10000101), .in_free(out_router134), .in_r1R(l_min[141]), .in_r2R(l_max[142]), .in_r1L(r_min[125]), .in_r2L(r_max[124]), .out_r1R(r_min[133]), .out_r2R(r_max[133]), .out_r1L(l_min[133]), .out_r2L(l_max[133]), .out_data(out_data[133]));
	apo_router_144_nodes r135 (.clk(clk), .router_name(8'b10000110), .in_free(out_router135), .in_r1R(l_min[142]), .in_r2R(l_max[143]), .in_r1L(r_min[126]), .in_r2L(r_max[125]), .out_r1R(r_min[134]), .out_r2R(r_max[134]), .out_r1L(l_min[134]), .out_r2L(l_max[134]), .out_data(out_data[134]));
	apo_router_144_nodes r136 (.clk(clk), .router_name(8'b10000111), .in_free(out_router136), .in_r1R(l_min[143]), .in_r2R(l_max[0]), .in_r1L(r_min[127]), .in_r2L(r_max[126]), .out_r1R(r_min[135]), .out_r2R(r_max[135]), .out_r1L(l_min[135]), .out_r2L(l_max[135]), .out_data(out_data[135]));
	apo_router_144_nodes r137 (.clk(clk), .router_name(8'b10001000), .in_free(out_router137), .in_r1R(l_min[0]), .in_r2R(l_max[1]), .in_r1L(r_min[128]), .in_r2L(r_max[127]), .out_r1R(r_min[136]), .out_r2R(r_max[136]), .out_r1L(l_min[136]), .out_r2L(l_max[136]), .out_data(out_data[136]));
	apo_router_144_nodes r138 (.clk(clk), .router_name(8'b10001001), .in_free(out_router138), .in_r1R(l_min[1]), .in_r2R(l_max[2]), .in_r1L(r_min[129]), .in_r2L(r_max[128]), .out_r1R(r_min[137]), .out_r2R(r_max[137]), .out_r1L(l_min[137]), .out_r2L(l_max[137]), .out_data(out_data[137]));
	apo_router_144_nodes r139 (.clk(clk), .router_name(8'b10001010), .in_free(out_router139), .in_r1R(l_min[2]), .in_r2R(l_max[3]), .in_r1L(r_min[130]), .in_r2L(r_max[129]), .out_r1R(r_min[138]), .out_r2R(r_max[138]), .out_r1L(l_min[138]), .out_r2L(l_max[138]), .out_data(out_data[138]));
	apo_router_144_nodes r140 (.clk(clk), .router_name(8'b10001011), .in_free(out_router140), .in_r1R(l_min[3]), .in_r2R(l_max[4]), .in_r1L(r_min[131]), .in_r2L(r_max[130]), .out_r1R(r_min[139]), .out_r2R(r_max[139]), .out_r1L(l_min[139]), .out_r2L(l_max[139]), .out_data(out_data[139]));
	apo_router_144_nodes r141 (.clk(clk), .router_name(8'b10001100), .in_free(out_router141), .in_r1R(l_min[4]), .in_r2R(l_max[5]), .in_r1L(r_min[132]), .in_r2L(r_max[131]), .out_r1R(r_min[140]), .out_r2R(r_max[140]), .out_r1L(l_min[140]), .out_r2L(l_max[140]), .out_data(out_data[140]));
	apo_router_144_nodes r142 (.clk(clk), .router_name(8'b10001101), .in_free(out_router142), .in_r1R(l_min[5]), .in_r2R(l_max[6]), .in_r1L(r_min[133]), .in_r2L(r_max[132]), .out_r1R(r_min[141]), .out_r2R(r_max[141]), .out_r1L(l_min[141]), .out_r2L(l_max[141]), .out_data(out_data[141]));
	apo_router_144_nodes r143 (.clk(clk), .router_name(8'b10001110), .in_free(out_router143), .in_r1R(l_min[6]), .in_r2R(l_max[7]), .in_r1L(r_min[134]), .in_r2L(r_max[133]), .out_r1R(r_min[142]), .out_r2R(r_max[142]), .out_r1L(l_min[142]), .out_r2L(l_max[142]), .out_data(out_data[142]));
	apo_router_144_nodes r144 (.clk(clk), .router_name(8'b10001111), .in_free(out_router144), .in_r1R(l_min[7]), .in_r2R(l_max[8]), .in_r1L(r_min[135]), .in_r2L(r_max[134]), .out_r1R(r_min[143]), .out_r2R(r_max[143]), .out_r1L(l_min[143]), .out_r2L(l_max[143]), .out_data(out_data[143]));

endmodule

